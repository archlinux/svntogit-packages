### start sv
DICT sv SE sv_SE
HYPH sv SE hyph_sv_SE
### end sv